module pixel_gen
(
input wire rst,
input wire [9:0]x_pxl,y_pxl,
output wire [11:0]rgb
);
//RGB12[(x_pxl*4'd3)+(12'd354*y_pxl)],RGB12[(x_pxl*4'd3)+(12'd354*y_pxl)+4'd1],RGB12[(x_pxl*4'd3)+(12'd354*y_pxl)+4'd2]
//101952'h...  {4'b0000,{4{1'b1}},4'b0000}
reg  [3:0] RGB12[0:25487]='{4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'h2,4'h2,4'h2,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h1,4'h1,4'h1,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'h1,4'h1,4'h1,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h0,4'h0,4'h0,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h6,4'h6,4'h6,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h1,4'h1,4'h1,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h0,4'h0,4'h0,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'hE,4'hE,4'hE,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h2,4'h2,4'h2,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'h0,4'h0,4'h0,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h0,4'h0,4'h0,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h1,4'h1,4'h1,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'h0,4'h0,4'h0,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h1,4'h1,4'h1,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'hB,4'hB,4'hB,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h1,4'h1,4'h1,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'h1,4'h1,4'h1,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h2,4'h2,4'h2,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h4,4'h4,4'h4,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h5,4'h5,4'h5,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h8,4'h8,4'h8,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hA,4'hA,4'hA,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h8,4'h8,4'h8,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'hA,4'hA,4'hA,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'hB,4'hB,4'hB,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h6,4'h6,4'h6,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'hA,4'hA,4'hA,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h9,4'h9,4'h9,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hB,4'hB,4'hB,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'h6,4'h6,4'h6,4'h0,4'h0,4'h0,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h6,4'h6,4'h6,4'hA,4'hA,4'hA,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h8,4'h8,4'h8,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h3,4'h3,4'h3,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hE,4'hE,4'hE,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h4,4'h4,4'h4,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hD,4'hD,4'hD,4'h7,4'h7,4'h7,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hE,4'hE,4'hE,4'hC,4'hC,4'hC,4'hF,4'hF,4'hF,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h9,4'h9,4'h9,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h6,4'h6,4'h6,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h5,4'h5,4'h5,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hC,4'hC,4'hC,4'h9,4'h9,4'h9,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h0,4'h0,4'h0,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h5,4'h5,4'h5,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'h0,4'h0,4'h0,4'h7,4'h7,4'h7,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h6,4'h6,4'h6,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h5,4'h5,4'h5,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h2,4'h2,4'h2,4'h2,4'h2,4'h2,4'h3,4'h3,4'h3,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'h0,4'h0,4'h0,4'h3,4'h3,4'h3,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h4,4'h4,4'h4,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h4,4'h4,4'h4,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h5,4'h5,4'h5,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h3,4'h2,4'h2,4'h2,4'h0,4'h0,4'h0,4'h4,4'h4,4'h4,4'h3,4'h3,4'h3,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hD,4'hD,4'hD,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h3,4'h3,4'h3,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h1,4'h0,4'h0,4'h0,4'h0,4'h0,4'h0,4'h5,4'h5,4'h5,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h6,4'h6,4'h6,4'h5,4'h5,4'h5,4'h4,4'h4,4'h4,4'h4,4'h4,4'h4,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h9,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'h8,4'h8,4'h8,4'h5,4'h5,4'h5,4'h2,4'h2,4'h2,4'h1,4'h1,4'h1,4'h5,4'h5,4'h5,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hE,4'hE,4'hE,4'hB,4'hB,4'hB,4'h8,4'h8,4'h8,4'h6,4'h6,4'h6,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hB,4'hB,4'hB,4'h9,4'h9,4'h9,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h8,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hC,4'hC,4'hC,4'hA,4'hA,4'hA,4'h7,4'h7,4'h7,4'h6,4'h6,4'h6,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h7,4'h8,4'h8,4'h8,4'h9,4'h9,4'h9,4'hB,4'hB,4'hB,4'hE,4'hE,4'hE,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hD,4'hD,4'hD,4'hC,4'hC,4'hC,4'hB,4'hB,4'hB,4'hA,4'hA,4'hA,4'hB,4'hB,4'hB,4'hC,4'hC,4'hC,4'hD,4'hD,4'hD,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF,4'hF};
//118x72 del_orean.png   
assign rgb = (x_pxl == 10'b1111111111 || y_pxl == 10'b1111111111) ? {24{1'b0}} :
				 ((x_pxl<=12'd117 && y_pxl<=16'd71 ) ? {RGB12[(x_pxl*12'd3)+(16'd354*y_pxl)], RGB12[(x_pxl*12'd3)+(16'd354*y_pxl)+16'd1], RGB12[(x_pxl*12'd3)+(16'd354*y_pxl)+16'd2]}:
				 12'h999);

endmodule